package memory_pkg;
	
	import uvm_pkg::*;
	import apb_master_pkg::*;
	import apb_slave_pkg::*;
	import apb_common_pkg::*;

        `include "memory_defines.svh"
	`include "uvm_macros.svh"
	`include "apb_base_seq_item.svh"
	`include "memory_sequencer.svh"
	`include "memory_driver.svh"
	`include "memory_agent.svh"
	`include "memory_env.svh"
	`include "memory_test.svh"


endpackage
