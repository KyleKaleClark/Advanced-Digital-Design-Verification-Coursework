module even_odd
(
	input 	clk, reset, w_en, r_en,
	input 	[7:0] d_in,
	output 	[7:0] d_out
);



endmodule
