a21164_asu@nc-asu6-l01.apporto.com.62288:1751758680