module fifo_tb();
	initial begin
		$display("hello world");
	end
endmodule
