`ifndef MEM_DEFINES
`define MEM_DEFINES

`define AWIDTH 10
`define DWIDTH 8
`define MAT_MUL_SIZE 4

typedef enum {READ, WRITE} mem_op_t;		

`endif
