package memory_pkg;
	
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "memory_interface.svh"
	`include "memory_driver.svh"
	`include "memory_agent.svh"
	`include "memory_sequencer.svh"
	`include "memory_env.svh"
	`include "memory_test.svh"

endpackage
